module top_module (
    input a,
    input b,
    input c,
    input d,
    output q );//

    assign q =~(a | b)?1'b0:(c|d); 

endmodule
